module adder (
    input [7:0] In,
    Output [7:0] Out
);

assign Out = In + 1 ;
    
endmodule